
`include "./../sysconfig.v"

/**
* 取指模块
*/
module fetch (
    //指令地址
    input wire [`XLEN-1:0] inst_addr,
    //指令内容
    output wire [`INST_LEN-1:0] inst_data
);


endmodule
