`include "./../sysconfig.v"


module clint (
    input clk,
    input rst
);

endmodule
