// lab01 开关实验
module lab01switch(
    input a,
    input b,
    output f
  );
  assign f = a ^ b;

endmodule
