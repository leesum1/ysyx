module writeback ();

endmodule
